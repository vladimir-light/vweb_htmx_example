module controllers
import vweb

struct IndexController {
	vweb.Context
}
